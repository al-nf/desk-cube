module led(
    output wire led0_r
);

    assign led0_r = 1'b1;

endmodule